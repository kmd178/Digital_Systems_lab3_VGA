`timescale 1ns / 1ps

module vga_testImage_BRAM_initialization_BLUE(
    );


endmodule
