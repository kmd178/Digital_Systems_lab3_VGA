`timescale 1ns / 1ps
module vga_controller(
input reset, 
input clk, 
output VGA_RED,
output VGA_GREEN,
output VGA_BLUE,
output VGA_HSYNC, 
output VGA_VSYNC);

endmodule
