
module vga_testImage_BRAM_initialization_GREEN(
    );


endmodule
